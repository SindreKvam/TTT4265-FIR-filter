library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ieee_proposed;
use ieee_proposed.fixed_float_types.all; -- ieee_proposed for VHDL-93 version
use ieee_proposed.fixed_pkg.all; -- ieee_proposed for compatibility version

entity fir is
    generic (
        FIR_LENGTH : integer
    );
    port (
        clk : in std_logic;
        rst_n : in std_logic;

        prev_ready : out std_logic;
        prev_valid : in std_logic;
        data_in : in std_logic_vector(0 downto 0);

        next_ready : in std_logic;
        next_valid : out std_logic;
        data_out : out sfixed(0 downto -23)
    );
end fir;

architecture rtl of fir is

    type T_STATE is (IDLE, SHIFT_DATA_IN, CALCULATE, HOLD_DATA_OUT);
    signal state : T_STATE := IDLE;

    type T_DATA is array(0 to FIR_LENGTH - 1) of std_logic_vector(0 downto 0); -- 1 bit
    signal delay_line : T_DATA := (others => (others => '0'));

    type T_COEFF is array(0 to FIR_LENGTH - 1) of sfixed(0 downto -21); -- 22 bit
    signal coeff : T_COEFF :=  ("11"&x"FFD26", "11"&x"FF7D8", "11"&x"FF3AF", "11"&x"FF141", "11"&x"FF0E6", "11"&x"FF2AB", "11"&x"FF651", "11"&x"FFB54", "00"&x"00100", "00"&x"00689", "00"&x"00B27", "00"&x"00E34", "00"&x"00F42", "00"&x"00E29", "00"&x"00B13", "00"&x"0066D", 
                                "00"&x"000DE", "11"&x"FFB2F", "11"&x"FF62D", "11"&x"FF28C", "11"&x"FF0D0", "11"&x"FF136", "11"&x"FF3B1", "11"&x"FF7E8", "11"&x"FFD43", "00"&x"00302", "00"&x"00855", "00"&x"00C7C", "00"&x"00EE2", "00"&x"00F30", "00"&x"00D5B", "00"&x"009A4", 
                                "00"&x"00491", "11"&x"FFED9", "11"&x"FF949", "11"&x"FF4AB", "11"&x"FF1A4", "11"&x"FF0A2", "11"&x"FF1C9", "11"&x"FF4F1", "11"&x"FF9A8", "11"&x"FFF44", "00"&x"004FB", "00"&x"009FF", "00"&x"00D9C", "00"&x"00F4F", "00"&x"00EDA", "00"&x"00C4F", 
                                "00"&x"00807", "00"&x"0029D", "11"&x"FFCD4", "11"&x"FF77D", "11"&x"FF358", "11"&x"FF0FA", "11"&x"FF0B9", "11"&x"FF29E", "11"&x"FF666", "11"&x"FFB88", "00"&x"0014C", "00"&x"006E2", "00"&x"00B81", "00"&x"00E81", "00"&x"00F77", "00"&x"00E40", 
                                "00"&x"00B08", "00"&x"00641", "00"&x"00098", "11"&x"FFAD9", "11"&x"FF5D3", "11"&x"FF23B", "11"&x"FF092", "11"&x"FF115", "11"&x"FF3B2", "11"&x"FF80A", "11"&x"FFD82", "00"&x"00354", "00"&x"008AF", "00"&x"00CD1", "00"&x"00F27", "00"&x"00F5A", 
                                "00"&x"00D65", "00"&x"0098C", "00"&x"0045B", "11"&x"FFE8C", "11"&x"FF8F1", "11"&x"FF453", "11"&x"FF159", "11"&x"FF06F", "11"&x"FF1B6", "11"&x"FF4FF", "11"&x"FF9D6", "11"&x"FFF8B", "00"&x"00551", "00"&x"00A58", "00"&x"00DEB", "00"&x"00F89", 
                                "00"&x"00EF8", "00"&x"00C4A", "00"&x"007E2", "00"&x"0025D", "11"&x"FFC82", "11"&x"FF724", "11"&x"FF305", "11"&x"FF0B8", "11"&x"FF092", "11"&x"FF298", "11"&x"FF681", "11"&x"FFBC1", "00"&x"0019A", "00"&x"0073A", "00"&x"00BD6", "00"&x"00EC9", 
                                "00"&x"00FA7", "00"&x"00E50", "00"&x"00AF6", "00"&x"00611", "00"&x"00050", "11"&x"FFA83", "11"&x"FF57C", "11"&x"FF1EE", "11"&x"FF05B", "11"&x"FF0FB", "11"&x"FF3B9", "11"&x"FF831", "11"&x"FFDC3", "00"&x"003A6", "00"&x"00907", "00"&x"00D22", 
                                "00"&x"00F65", "00"&x"00F7D", "00"&x"00D67", "00"&x"0096E", "00"&x"00421", "11"&x"FFE3E", "11"&x"FF89A", "11"&x"FF3FF", "11"&x"FF115", "11"&x"FF044", "11"&x"FF1A9", "11"&x"FF514", "11"&x"FFA08", "11"&x"FFFD4", "00"&x"005A6", "00"&x"00AAE", 
                                "00"&x"00E35", "00"&x"00FBD", "00"&x"00F0E", "00"&x"00C40", "00"&x"007B8", "00"&x"0021A", "11"&x"FFC2F", "11"&x"FF6CD", "11"&x"FF2B6", "11"&x"FF07D", "11"&x"FF073", "11"&x"FF299", "11"&x"FF6A2", "11"&x"FFBFD", "00"&x"001E9", "00"&x"00790", 
                                "00"&x"00C28", "00"&x"00F0A", "00"&x"00FCF", "00"&x"00E59", "00"&x"00ADF", "00"&x"005DD", "00"&x"00006", "11"&x"FFA2E", "11"&x"FF527", "11"&x"FF1A7", "11"&x"FF02B", "11"&x"FF0E9", "11"&x"FF3C7", "11"&x"FF85D", "11"&x"FFE07", "00"&x"003F9", 
                                "00"&x"0095C", "00"&x"00D6E", "00"&x"00F9D", "00"&x"00F99", "00"&x"00D63", "00"&x"0094B", "00"&x"003E3", "11"&x"FFDEF", "11"&x"FF844", "11"&x"FF3B0", "11"&x"FF0D6", "11"&x"FF01F", "11"&x"FF1A4", "11"&x"FF52E", "11"&x"FFA3E", "00"&x"0001E", 
                                "00"&x"005FB", "00"&x"00B00", "00"&x"00E7A", "00"&x"00FEA", "00"&x"00F1D", "00"&x"00C2F", "00"&x"0078A", "00"&x"001D5", "11"&x"FFBDD", "11"&x"FF67A", "11"&x"FF26D", "11"&x"FF049", "11"&x"FF05B", "11"&x"FF2A0", "11"&x"FF6C8", "11"&x"FFC3C", 
                                "00"&x"00238", "00"&x"007E5", "00"&x"00C75", "00"&x"00F46", "00"&x"00FF0", "00"&x"00E5C", "00"&x"00AC2", "00"&x"005A4", "11"&x"FFFBB", "11"&x"FF9DB", "11"&x"FF4D7", "11"&x"FF165", "11"&x"FF001", "11"&x"FF0DD", "11"&x"FF3DB", "11"&x"FF88E", 
                                "11"&x"FFE4E", "00"&x"0044B", "00"&x"009AE", "00"&x"00DB5", "00"&x"00FCE", "00"&x"00FAE", "00"&x"00D58", "00"&x"00922", "00"&x"003A2", "11"&x"FFD9F", "11"&x"FF7F1", "11"&x"FF365", "11"&x"FF09E", "11"&x"FF002", "11"&x"FF1A5", "11"&x"FF54E", 
                                "11"&x"FFA78", "00"&x"0006A", "00"&x"0064E", "00"&x"00B4E", "00"&x"00EB8", "00"&x"01010", "00"&x"00F25", "00"&x"00C18", "00"&x"00757", "00"&x"0018D", "11"&x"FFB8B", "11"&x"FF629", "11"&x"FF229", "11"&x"FF01B", "11"&x"FF04A", "11"&x"FF2AE", 
                                "11"&x"FF6F3", "11"&x"FFC7E", "00"&x"00288", "00"&x"00837", "00"&x"00CBE", "00"&x"00F7B", "00"&x"01009", "00"&x"00E57", "00"&x"00A9F", "00"&x"00568", "11"&x"FFF6E", "11"&x"FF988", "11"&x"FF48B", "11"&x"FF12A", "11"&x"FEFDF", "11"&x"FF0D9", 
                                "11"&x"FF3F5", "11"&x"FF8C3", "11"&x"FFE96", "00"&x"0049D", "00"&x"009FD", "00"&x"00DF6", "00"&x"00FF8", "00"&x"00FBB", "00"&x"00D47", "00"&x"008F4", "00"&x"0035F", "11"&x"FFD4F", "11"&x"FF7A0", "11"&x"FF31F", "11"&x"FF06C", "11"&x"FEFEB", 
                                "11"&x"FF1AD", "11"&x"FF574", "11"&x"FFAB6", "00"&x"000B7", "00"&x"0069F", "00"&x"00B99", "00"&x"00EF1", "00"&x"0102E", "00"&x"00F25", "00"&x"00BFA", "00"&x"00720", "00"&x"00144", "11"&x"FFB3A", "11"&x"FF5DC", "11"&x"FF1EA", "11"&x"FEFF4", 
                                "11"&x"FF040", "11"&x"FF2C3", "11"&x"FF723", "11"&x"FFCC3", "00"&x"002D8", "00"&x"00886", "00"&x"00D02", "00"&x"00FA9", "00"&x"0101C", "00"&x"00E4B", "00"&x"00A76", "00"&x"00529", "11"&x"FFF21", "11"&x"FF938", "11"&x"FF443", "11"&x"FF0F5", 
                                "11"&x"FEFC4", "11"&x"FF0DC", "11"&x"FF416", "11"&x"FF8FD", "11"&x"FFEE0", "00"&x"004ED", "00"&x"00A48", "00"&x"00E32", "00"&x"0101B", "00"&x"00FC1", "00"&x"00D2F", "00"&x"008C2", "00"&x"00319", "11"&x"FFD00", "11"&x"FF753", "11"&x"FF2DE", 
                                "11"&x"FF042", "11"&x"FEFDC", "11"&x"FF1BD", "11"&x"FF59F", "11"&x"FFAF7", "00"&x"00105", "00"&x"006EE", "00"&x"00BDE", "00"&x"00F23", "00"&x"01046", "00"&x"00F1F", "00"&x"00BD7", "00"&x"006E4", "00"&x"000F9", "11"&x"FFAEA", "11"&x"FF592", 
                                "11"&x"FF1B2", "11"&x"FEFD5", "11"&x"FF03E", "11"&x"FF2DE", "11"&x"FF758", "11"&x"FFD0A", "00"&x"00327", "00"&x"008D2", "00"&x"00D40", "00"&x"00FD0", "00"&x"01027", "00"&x"00E38", "00"&x"00A48", "00"&x"004E6", "11"&x"FFED3", "11"&x"FF8EA", 
                                "11"&x"FF400", "11"&x"FF0C6", "11"&x"FEFB0", "11"&x"FF0E6", "11"&x"FF43C", "11"&x"FF93A", "11"&x"FFF2C", "00"&x"0053C", "00"&x"00A90", "00"&x"00E67", "00"&x"01038", "00"&x"00FC0", "00"&x"00D11", "00"&x"0088B", "00"&x"002D1", "11"&x"FFCB1", 
                                "11"&x"FF708", "11"&x"FF2A2", "11"&x"FF01D", "11"&x"FEFD5", "11"&x"FF1D3", "11"&x"FF5CF", "11"&x"FFB3B", "00"&x"00153", "00"&x"0073B", "00"&x"00C1F", "00"&x"00F4E", "00"&x"01056", "00"&x"00F11", "00"&x"00BAE", "00"&x"006A5", "00"&x"000AD", 
                                "11"&x"FFA9C", "11"&x"FF54D", "11"&x"FF180", "11"&x"FEFBC", "11"&x"FF043", "11"&x"FF300", "11"&x"FF792", "11"&x"FFD53", "00"&x"00375", "00"&x"0091B", "00"&x"00D79", "00"&x"00FF1", "00"&x"0102B", "00"&x"00E1F", "00"&x"00A15", "00"&x"004A1", 
                                "11"&x"FFE85", "11"&x"FF89F", "11"&x"FF3C2", "11"&x"FF09E", "11"&x"FEFA4", "11"&x"FF0F7", "11"&x"FF468", "11"&x"FF97B", "11"&x"FFF78", "00"&x"00589", "00"&x"00AD3", "00"&x"00E96", "00"&x"0104C", "00"&x"00FB7", "00"&x"00CEC", "00"&x"0084F", 
                                "00"&x"00286", "11"&x"FFC63", "11"&x"FF6C1", "11"&x"FF26C", "11"&x"FF000", "11"&x"FEFD5", "11"&x"FF1F0", "11"&x"FF605", "11"&x"FFB82", "00"&x"001A1", "00"&x"00785", "00"&x"00C5A", "00"&x"00F73", "00"&x"0105F", "00"&x"00EFD", "00"&x"00B7F", 
                                "00"&x"00663", "00"&x"00060", "11"&x"FFA50", "11"&x"FF50D", "11"&x"FF154", "11"&x"FEFAB", "11"&x"FF04F", "11"&x"FF328", "11"&x"FF7CF", "11"&x"FFD9E", "00"&x"003C3", "00"&x"00960", "00"&x"00DAB", "00"&x"0100A", "00"&x"01027", "00"&x"00DFF", 
                                "00"&x"009DD", "00"&x"00459", "11"&x"FFE37", "11"&x"FF856", "11"&x"FF389", "11"&x"FF07C", "11"&x"FEF9F", "11"&x"FF10F", "11"&x"FF49A", "11"&x"FF9BF", "11"&x"FFFC5", "00"&x"005D4", "00"&x"00B11", "00"&x"00EBF", "00"&x"0105A", "00"&x"00FA8", 
                                "00"&x"00CC1", "00"&x"0080F", "00"&x"0023B", "11"&x"FFC16", "11"&x"FF67E", "11"&x"FF23D", "11"&x"FEFEB", "11"&x"FEFDC", "11"&x"FF213", "11"&x"FF63F", "11"&x"FFBCB", "00"&x"001EE", "00"&x"007CC", "00"&x"00C91", "00"&x"00F91", "00"&x"01060", 
                                "00"&x"00EE1", "00"&x"00B4A", "00"&x"0061D", "00"&x"00013", "11"&x"FFA06", "11"&x"FF4D1", "11"&x"FF12E", "11"&x"FEFA1", "11"&x"FF062", "11"&x"FF355", "11"&x"FF811", "11"&x"FFDEA", "00"&x"0040F", "00"&x"009A1", "00"&x"00DD8", "00"&x"0101D", 
                                "00"&x"0101D", "00"&x"00DD8", "00"&x"009A1", "00"&x"0040F", "11"&x"FFDEA", "11"&x"FF811", "11"&x"FF355", "11"&x"FF062", "11"&x"FEFA1", "11"&x"FF12E", "11"&x"FF4D1", "11"&x"FFA06", "00"&x"00013", "00"&x"0061D", "00"&x"00B4A", "00"&x"00EE1", 
                                "00"&x"01060", "00"&x"00F91", "00"&x"00C91", "00"&x"007CC", "00"&x"001EE", "11"&x"FFBCB", "11"&x"FF63F", "11"&x"FF213", "11"&x"FEFDC", "11"&x"FEFEB", "11"&x"FF23D", "11"&x"FF67E", "11"&x"FFC16", "00"&x"0023B", "00"&x"0080F", "00"&x"00CC1", 
                                "00"&x"00FA8", "00"&x"0105A", "00"&x"00EBF", "00"&x"00B11", "00"&x"005D4", "11"&x"FFFC5", "11"&x"FF9BF", "11"&x"FF49A", "11"&x"FF10F", "11"&x"FEF9F", "11"&x"FF07C", "11"&x"FF389", "11"&x"FF856", "11"&x"FFE37", "00"&x"00459", "00"&x"009DD", 
                                "00"&x"00DFF", "00"&x"01027", "00"&x"0100A", "00"&x"00DAB", "00"&x"00960", "00"&x"003C3", "11"&x"FFD9E", "11"&x"FF7CF", "11"&x"FF328", "11"&x"FF04F", "11"&x"FEFAB", "11"&x"FF154", "11"&x"FF50D", "11"&x"FFA50", "00"&x"00060", "00"&x"00663", 
                                "00"&x"00B7F", "00"&x"00EFD", "00"&x"0105F", "00"&x"00F73", "00"&x"00C5A", "00"&x"00785", "00"&x"001A1", "11"&x"FFB82", "11"&x"FF605", "11"&x"FF1F0", "11"&x"FEFD5", "11"&x"FF000", "11"&x"FF26C", "11"&x"FF6C1", "11"&x"FFC63", "00"&x"00286", 
                                "00"&x"0084F", "00"&x"00CEC", "00"&x"00FB7", "00"&x"0104C", "00"&x"00E96", "00"&x"00AD3", "00"&x"00589", "11"&x"FFF78", "11"&x"FF97B", "11"&x"FF468", "11"&x"FF0F7", "11"&x"FEFA4", "11"&x"FF09E", "11"&x"FF3C2", "11"&x"FF89F", "11"&x"FFE85", 
                                "00"&x"004A1", "00"&x"00A15", "00"&x"00E1F", "00"&x"0102B", "00"&x"00FF1", "00"&x"00D79", "00"&x"0091B", "00"&x"00375", "11"&x"FFD53", "11"&x"FF792", "11"&x"FF300", "11"&x"FF043", "11"&x"FEFBC", "11"&x"FF180", "11"&x"FF54D", "11"&x"FFA9C", 
                                "00"&x"000AD", "00"&x"006A5", "00"&x"00BAE", "00"&x"00F11", "00"&x"01056", "00"&x"00F4E", "00"&x"00C1F", "00"&x"0073B", "00"&x"00153", "11"&x"FFB3B", "11"&x"FF5CF", "11"&x"FF1D3", "11"&x"FEFD5", "11"&x"FF01D", "11"&x"FF2A2", "11"&x"FF708", 
                                "11"&x"FFCB1", "00"&x"002D1", "00"&x"0088B", "00"&x"00D11", "00"&x"00FC0", "00"&x"01038", "00"&x"00E67", "00"&x"00A90", "00"&x"0053C", "11"&x"FFF2C", "11"&x"FF93A", "11"&x"FF43C", "11"&x"FF0E6", "11"&x"FEFB0", "11"&x"FF0C6", "11"&x"FF400", 
                                "11"&x"FF8EA", "11"&x"FFED3", "00"&x"004E6", "00"&x"00A48", "00"&x"00E38", "00"&x"01027", "00"&x"00FD0", "00"&x"00D40", "00"&x"008D2", "00"&x"00327", "11"&x"FFD0A", "11"&x"FF758", "11"&x"FF2DE", "11"&x"FF03E", "11"&x"FEFD5", "11"&x"FF1B2", 
                                "11"&x"FF592", "11"&x"FFAEA", "00"&x"000F9", "00"&x"006E4", "00"&x"00BD7", "00"&x"00F1F", "00"&x"01046", "00"&x"00F23", "00"&x"00BDE", "00"&x"006EE", "00"&x"00105", "11"&x"FFAF7", "11"&x"FF59F", "11"&x"FF1BD", "11"&x"FEFDC", "11"&x"FF042", 
                                "11"&x"FF2DE", "11"&x"FF753", "11"&x"FFD00", "00"&x"00319", "00"&x"008C2", "00"&x"00D2F", "00"&x"00FC1", "00"&x"0101B", "00"&x"00E32", "00"&x"00A48", "00"&x"004ED", "11"&x"FFEE0", "11"&x"FF8FD", "11"&x"FF416", "11"&x"FF0DC", "11"&x"FEFC4", 
                                "11"&x"FF0F5", "11"&x"FF443", "11"&x"FF938", "11"&x"FFF21", "00"&x"00529", "00"&x"00A76", "00"&x"00E4B", "00"&x"0101C", "00"&x"00FA9", "00"&x"00D02", "00"&x"00886", "00"&x"002D8", "11"&x"FFCC3", "11"&x"FF723", "11"&x"FF2C3", "11"&x"FF040", 
                                "11"&x"FEFF4", "11"&x"FF1EA", "11"&x"FF5DC", "11"&x"FFB3A", "00"&x"00144", "00"&x"00720", "00"&x"00BFA", "00"&x"00F25", "00"&x"0102E", "00"&x"00EF1", "00"&x"00B99", "00"&x"0069F", "00"&x"000B7", "11"&x"FFAB6", "11"&x"FF574", "11"&x"FF1AD", 
                                "11"&x"FEFEB", "11"&x"FF06C", "11"&x"FF31F", "11"&x"FF7A0", "11"&x"FFD4F", "00"&x"0035F", "00"&x"008F4", "00"&x"00D47", "00"&x"00FBB", "00"&x"00FF8", "00"&x"00DF6", "00"&x"009FD", "00"&x"0049D", "11"&x"FFE96", "11"&x"FF8C3", "11"&x"FF3F5", 
                                "11"&x"FF0D9", "11"&x"FEFDF", "11"&x"FF12A", "11"&x"FF48B", "11"&x"FF988", "11"&x"FFF6E", "00"&x"00568", "00"&x"00A9F", "00"&x"00E57", "00"&x"01009", "00"&x"00F7B", "00"&x"00CBE", "00"&x"00837", "00"&x"00288", "11"&x"FFC7E", "11"&x"FF6F3", 
                                "11"&x"FF2AE", "11"&x"FF04A", "11"&x"FF01B", "11"&x"FF229", "11"&x"FF629", "11"&x"FFB8B", "00"&x"0018D", "00"&x"00757", "00"&x"00C18", "00"&x"00F25", "00"&x"01010", "00"&x"00EB8", "00"&x"00B4E", "00"&x"0064E", "00"&x"0006A", "11"&x"FFA78", 
                                "11"&x"FF54E", "11"&x"FF1A5", "11"&x"FF002", "11"&x"FF09E", "11"&x"FF365", "11"&x"FF7F1", "11"&x"FFD9F", "00"&x"003A2", "00"&x"00922", "00"&x"00D58", "00"&x"00FAE", "00"&x"00FCE", "00"&x"00DB5", "00"&x"009AE", "00"&x"0044B", "11"&x"FFE4E", 
                                "11"&x"FF88E", "11"&x"FF3DB", "11"&x"FF0DD", "11"&x"FF001", "11"&x"FF165", "11"&x"FF4D7", "11"&x"FF9DB", "11"&x"FFFBB", "00"&x"005A4", "00"&x"00AC2", "00"&x"00E5C", "00"&x"00FF0", "00"&x"00F46", "00"&x"00C75", "00"&x"007E5", "00"&x"00238", 
                                "11"&x"FFC3C", "11"&x"FF6C8", "11"&x"FF2A0", "11"&x"FF05B", "11"&x"FF049", "11"&x"FF26D", "11"&x"FF67A", "11"&x"FFBDD", "00"&x"001D5", "00"&x"0078A", "00"&x"00C2F", "00"&x"00F1D", "00"&x"00FEA", "00"&x"00E7A", "00"&x"00B00", "00"&x"005FB", 
                                "00"&x"0001E", "11"&x"FFA3E", "11"&x"FF52E", "11"&x"FF1A4", "11"&x"FF01F", "11"&x"FF0D6", "11"&x"FF3B0", "11"&x"FF844", "11"&x"FFDEF", "00"&x"003E3", "00"&x"0094B", "00"&x"00D63", "00"&x"00F99", "00"&x"00F9D", "00"&x"00D6E", "00"&x"0095C", 
                                "00"&x"003F9", "11"&x"FFE07", "11"&x"FF85D", "11"&x"FF3C7", "11"&x"FF0E9", "11"&x"FF02B", "11"&x"FF1A7", "11"&x"FF527", "11"&x"FFA2E", "00"&x"00006", "00"&x"005DD", "00"&x"00ADF", "00"&x"00E59", "00"&x"00FCF", "00"&x"00F0A", "00"&x"00C28", 
                                "00"&x"00790", "00"&x"001E9", "11"&x"FFBFD", "11"&x"FF6A2", "11"&x"FF299", "11"&x"FF073", "11"&x"FF07D", "11"&x"FF2B6", "11"&x"FF6CD", "11"&x"FFC2F", "00"&x"0021A", "00"&x"007B8", "00"&x"00C40", "00"&x"00F0E", "00"&x"00FBD", "00"&x"00E35", 
                                "00"&x"00AAE", "00"&x"005A6", "11"&x"FFFD4", "11"&x"FFA08", "11"&x"FF514", "11"&x"FF1A9", "11"&x"FF044", "11"&x"FF115", "11"&x"FF3FF", "11"&x"FF89A", "11"&x"FFE3E", "00"&x"00421", "00"&x"0096E", "00"&x"00D67", "00"&x"00F7D", "00"&x"00F65", 
                                "00"&x"00D22", "00"&x"00907", "00"&x"003A6", "11"&x"FFDC3", "11"&x"FF831", "11"&x"FF3B9", "11"&x"FF0FB", "11"&x"FF05B", "11"&x"FF1EE", "11"&x"FF57C", "11"&x"FFA83", "00"&x"00050", "00"&x"00611", "00"&x"00AF6", "00"&x"00E50", "00"&x"00FA7", 
                                "00"&x"00EC9", "00"&x"00BD6", "00"&x"0073A", "00"&x"0019A", "11"&x"FFBC1", "11"&x"FF681", "11"&x"FF298", "11"&x"FF092", "11"&x"FF0B8", "11"&x"FF305", "11"&x"FF724", "11"&x"FFC82", "00"&x"0025D", "00"&x"007E2", "00"&x"00C4A", "00"&x"00EF8", 
                                "00"&x"00F89", "00"&x"00DEB", "00"&x"00A58", "00"&x"00551", "11"&x"FFF8B", "11"&x"FF9D6", "11"&x"FF4FF", "11"&x"FF1B6", "11"&x"FF06F", "11"&x"FF159", "11"&x"FF453", "11"&x"FF8F1", "11"&x"FFE8C", "00"&x"0045B", "00"&x"0098C", "00"&x"00D65", 
                                "00"&x"00F5A", "00"&x"00F27", "00"&x"00CD1", "00"&x"008AF", "00"&x"00354", "11"&x"FFD82", "11"&x"FF80A", "11"&x"FF3B2", "11"&x"FF115", "11"&x"FF092", "11"&x"FF23B", "11"&x"FF5D3", "11"&x"FFAD9", "00"&x"00098", "00"&x"00641", "00"&x"00B08", 
                                "00"&x"00E40", "00"&x"00F77", "00"&x"00E81", "00"&x"00B81", "00"&x"006E2", "00"&x"0014C", "11"&x"FFB88", "11"&x"FF666", "11"&x"FF29E", "11"&x"FF0B9", "11"&x"FF0FA", "11"&x"FF358", "11"&x"FF77D", "11"&x"FFCD4", "00"&x"0029D", "00"&x"00807", 
                                "00"&x"00C4F", "00"&x"00EDA", "00"&x"00F4F", "00"&x"00D9C", "00"&x"009FF", "00"&x"004FB", "11"&x"FFF44", "11"&x"FF9A8", "11"&x"FF4F1", "11"&x"FF1C9", "11"&x"FF0A2", "11"&x"FF1A4", "11"&x"FF4AB", "11"&x"FF949", "11"&x"FFED9", "00"&x"00491", 
                                "00"&x"009A4", "00"&x"00D5B", "00"&x"00F30", "00"&x"00EE2", "00"&x"00C7C", "00"&x"00855", "00"&x"00302", "11"&x"FFD43", "11"&x"FF7E8", "11"&x"FF3B1", "11"&x"FF136", "11"&x"FF0D0", "11"&x"FF28C", "11"&x"FF62D", "11"&x"FFB2F", "00"&x"000DE", 
                                "00"&x"0066D", "00"&x"00B13", "00"&x"00E29", "00"&x"00F42", "00"&x"00E34", "00"&x"00B27", "00"&x"00689", "00"&x"00100", "11"&x"FFB54", "11"&x"FF651", "11"&x"FF2AB", "11"&x"FF0E6", "11"&x"FF141", "11"&x"FF3AF", "11"&x"FF7D8", "11"&x"FFD26");

    -- 24 bit accumulator
    signal accumulator : sfixed(0 downto -23) := (others => '0');
    -- 12 bit because max sum is 1286.28
    --signal accumulator : signed(23 downto 0) := (others => '0');
    signal sfixed_data_in : sfixed(0 downto 0) := (others => '0');

    signal tap_counter : unsigned(11 downto 0) := (others => '0');
    

begin

    FIR_PROC : process(clk)

        variable v_prev_ready : std_logic := '0';
        variable v_next_valid : std_logic := '0';
        variable v_index : integer range 0 to FIR_LENGTH * 2 - 1 := 0;
        variable v_coeff : sfixed(0 downto -21);
        variable v_delay_line : sfixed(0 downto 0);
        variable v_mult_result : sfixed(0 downto -21);

    begin
        
        if rising_edge(clk) then

            -- Default values
            v_prev_ready := '0';
            v_next_valid := '0';

            if rst_n = '0' then

                state <= IDLE;
                
            else
                
                case state is

                    -------------------------------
                    when IDLE =>
                        -------------------------------
                        v_prev_ready := '1';

                        if prev_valid = '1' then
                            state <= SHIFT_DATA_IN;
                        end if;

                    -------------------------------
                    when SHIFT_DATA_IN =>
                        -------------------------------
                        delay_line <= data_in & delay_line(delay_line'low to delay_line'high - 1);

                        -- Get accumulator ready
                        accumulator <=  (others => '0');
                        state <= CALCULATE;


                    -------------------------------
                    when CALCULATE =>
                        -------------------------------

                        v_index := to_integer(tap_counter);

                        v_coeff := coeff(v_index);
                        v_delay_line := to_sfixed(delay_line(v_index)(0 downto 0), v_delay_line);

                        v_mult_result := resize(v_coeff * v_delay_line , v_mult_result); -- * to_sfixed(-1, v_delay_line)

                        accumulator <= resize(accumulator + v_mult_result, accumulator);--fixed_saturate, fixed_round);

                        if (tap_counter < FIR_LENGTH - 1) then
                            tap_counter <= tap_counter + 1;
                        else
                            tap_counter <= (others => '0');
                            state <= HOLD_DATA_OUT;
                        end if;

                    -------------------------------
                    when HOLD_DATA_OUT =>
                        -------------------------------
                        v_next_valid := '1';

                        data_out <= accumulator;
                        
                        if next_ready = '1' then
                            state <= IDLE;
                        end if;

                    -------------------------------
                    when others => 
                        -------------------------------
                        state <= IDLE;

                end case;

            end if;

            prev_ready <= v_prev_ready;
            next_valid <= v_next_valid;

        end if;
        
    end process;

end architecture;