library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ieee_proposed;
use ieee_proposed.fixed_float_types.all; -- ieee_proposed for VHDL-93 version
use ieee_proposed.fixed_pkg.all; -- ieee_proposed for compatibility version

entity fir is
    generic (
        FIR_LENGTH : integer
    );
    port (
        clk : in std_logic;
        rst_n : in std_logic;

        prev_ready : out std_logic;
        prev_valid : in std_logic;
        data_in : in std_logic_vector(0 downto 0);

        next_ready : in std_logic;
        next_valid : out std_logic;
        data_out : out sfixed(0 downto -23)
    );
end fir;

architecture rtl of fir is

    type T_STATE is (IDLE, SHIFT_DATA_IN, CALCULATE, HOLD_DATA_OUT);
    signal state : T_STATE := IDLE;

    type T_DATA is array(0 to FIR_LENGTH - 1) of std_logic_vector(0 downto 0); -- 1 bit
    signal delay_line : T_DATA := (others => (others => '0'));

    type T_COEFF is array(0 to FIR_LENGTH - 1) of sfixed(0 downto -21); -- 22 bit
    signal coeff : T_COEFF :=  ("00"&x"005FC", "11"&x"FF272", "00"&x"00B44", "11"&x"FFF21", "11"&x"FF5F2", "00"&x"00D9D", "11"&x"FF8AF", "11"&x"FFBCD", "00"&x"00C8F", "11"&x"FF439", "00"&x"00280", "00"&x"00877", "11"&x"FF2CA", "00"&x"0085E", "00"&x"00272", "11"&x"FF4A1", 
                                "00"&x"00BFC", "11"&x"FFC0A", "11"&x"FF92E", "00"&x"00C8A", "11"&x"FF6D9", "11"&x"FFF37", "00"&x"00A03", "11"&x"FF418", "00"&x"00531", "00"&x"00527", "11"&x"FF45C", "00"&x"009A5", "11"&x"FFF41", "11"&x"FF772", "00"&x"00B8B", "11"&x"FF9D1", 
                                "11"&x"FFC77", "00"&x"00A8A", "11"&x"FF627", "00"&x"00216", "00"&x"00707", "11"&x"FF513", "00"&x"006E5", "00"&x"00201", "11"&x"FF6B5", "00"&x"009C1", "11"&x"FFCCA", "11"&x"FFA7E", "00"&x"00A14", "11"&x"FF8AD", "11"&x"FFF60", "00"&x"007F0", 
                                "11"&x"FF69B", "00"&x"00414", "00"&x"00407", "11"&x"FF6F4", "00"&x"00775", "11"&x"FFF6D", "11"&x"FF975", "00"&x"008C6", "11"&x"FFB53", "11"&x"FFD58", "00"&x"007DF", "11"&x"FF8B1", "00"&x"00189", "00"&x"00525", "11"&x"FF80E", "00"&x"004FA", 
                                "00"&x"00170", "11"&x"FF964", "00"&x"006E1", "11"&x"FFDC1", "11"&x"FFC2E", "00"&x"006EE", "11"&x"FFB02", "11"&x"FFF94", "00"&x"0054E", "11"&x"FF9C9", "00"&x"002AB", "00"&x"0029B", "11"&x"FFA36", "00"&x"004B7", "11"&x"FFFA4", "11"&x"FFBF8", 
                                "00"&x"00555", "11"&x"FFD33", "11"&x"FFE6E", "00"&x"00492", "11"&x"FFBD4", "00"&x"000DC", "00"&x"002D5", "11"&x"FFBB6", "00"&x"002A1", "00"&x"000BE", "11"&x"FFCAA", "00"&x"00363", "11"&x"FFEEC", "11"&x"FFE39", "00"&x"0031F", "11"&x"FFDD3", 
                                "11"&x"FFFD2", "00"&x"00223", "11"&x"FFD9A", "00"&x"000FB", "00"&x"000E8", "11"&x"FFE19", "00"&x"00172", "11"&x"FFFE6", "11"&x"FFEF3", "00"&x"00140", "11"&x"FFF6B", "11"&x"FFFB8", "00"&x"000AC", "11"&x"FFF85", "00"&x"00011", "00"&x"0001D", 
                                "00"&x"00000", "11"&x"FFFE1", "11"&x"FFFEE", "00"&x"0007C", "11"&x"FFF4F", "00"&x"00049", "00"&x"00099", "11"&x"FFEB4", "00"&x"00117", "00"&x"0001B", "11"&x"FFE7A", "00"&x"00201", "11"&x"FFF09", "11"&x"FFEF3", "00"&x"00292", "11"&x"FFDB1", 
                                "00"&x"00031", "00"&x"0025D", "11"&x"FFC95", "00"&x"001F3", "00"&x"00130", "11"&x"FFC3C", "00"&x"003B9", "11"&x"FFF2A", "11"&x"FFD08", "00"&x"004DB", "11"&x"FFCC5", "11"&x"FFF03", "00"&x"004CC", "11"&x"FFAB6", "00"&x"001D2", "00"&x"00345", 
                                "11"&x"FF9BC", "00"&x"004C1", "00"&x"0006C", "11"&x"FFA61", "00"&x"006EF", "11"&x"FFCDC", "11"&x"FFCC5", "00"&x"0078E", "11"&x"FF983", "00"&x"00084", "00"&x"00629", "11"&x"FF766", "00"&x"004C3", "00"&x"002D0", "11"&x"FF754", "00"&x"0085D", 
                                "11"&x"FFE2B", "11"&x"FF9A1", "00"&x"00A36", "11"&x"FF959", "11"&x"FFE00", "00"&x"00989", "11"&x"FF5AB", "00"&x"00380", "00"&x"00631", "11"&x"FF44E", "00"&x"008C2", "00"&x"000C4", "11"&x"FF5E9", "00"&x"00C4D", "11"&x"FFA7E", "11"&x"FFA65", 
                                "00"&x"00CF8", "11"&x"FF4FA", "00"&x"000DE", "00"&x"00A44", "11"&x"FF1CA", "00"&x"007CC", "00"&x"00491", "11"&x"FF208", "00"&x"00D5E", "11"&x"FFD18", "11"&x"FF5F9", "00"&x"00FF7", "11"&x"FF5AB", "11"&x"FFCEB", "00"&x"00E9D", "11"&x"FF045", 
                                "00"&x"0054D", "00"&x"00952", "11"&x"FEE80", "00"&x"00D07", "00"&x"00123", "11"&x"FF126", "00"&x"01203", "11"&x"FF7FA", "11"&x"FF7E0", "00"&x"012B7", "11"&x"FF02B", "00"&x"0013E", "00"&x"00E9E", "11"&x"FEBDC", "00"&x"00B01", "00"&x"0066C", 
                                "11"&x"FEC71", "00"&x"012A5", "11"&x"FFBF7", "11"&x"FF21F", "00"&x"01603", "11"&x"FF1CF", "11"&x"FFBC8", "00"&x"013F0", "11"&x"FEA9C", "00"&x"0072F", "00"&x"00C97", "11"&x"FE871", "00"&x"0117D", "00"&x"00185", "11"&x"FEC2F", "00"&x"017F6", 
                                "11"&x"FF55C", "11"&x"FF541", "00"&x"018AF", "11"&x"FEB2D", "00"&x"001A1", "00"&x"01320", "11"&x"FE5B8", "00"&x"00E53", "00"&x"00856", "11"&x"FE6AC", "00"&x"01816", "11"&x"FFACD", "11"&x"FEE28", "00"&x"01C3D", "11"&x"FEDD6", "11"&x"FFA9D", 
                                "00"&x"01968", "11"&x"FE4CF", "00"&x"0091D", "00"&x"00FF0", "11"&x"FE23D", "00"&x"0160C", "00"&x"001EA", "11"&x"FE71F", "00"&x"01E07", "11"&x"FF2B1", "11"&x"FF295", "00"&x"01EC2", "11"&x"FE61A", "00"&x"00206", "00"&x"017B2", "11"&x"FDF7F", 
                                "00"&x"011B0", "00"&x"00A47", "11"&x"FE0D6", "00"&x"01D96", "11"&x"FF9A0", "11"&x"FEA28", "00"&x"02284", "11"&x"FE9D6", "11"&x"FF970", "00"&x"01EE7", "11"&x"FDEFA", "00"&x"00B0D", "00"&x"0134C", "11"&x"FDC05", "00"&x"01A9E", "00"&x"0024E", 
                                "11"&x"FE20E", "00"&x"02417", "11"&x"FF007", "11"&x"FEFEC", "00"&x"024CF", "11"&x"FE10D", "00"&x"0026A", "00"&x"01C3E", "11"&x"FD950", "00"&x"01506", "00"&x"00C33", "11"&x"FDB0E", "00"&x"02308", "11"&x"FF876", "11"&x"FE634", "00"&x"028B6", 
                                "11"&x"FE5E4", "11"&x"FF847", "00"&x"02451", "11"&x"FD93C", "00"&x"00CF5", "00"&x"01699", "11"&x"FD5EA", "00"&x"01F18", "00"&x"002B1", "11"&x"FDD19", "00"&x"02A04", "11"&x"FED6D", "11"&x"FED53", "00"&x"02AB7", "11"&x"FDC20", "00"&x"002CC", 
                                "00"&x"020AB", "11"&x"FD34D", "00"&x"01844", "00"&x"00E11", "11"&x"FD573", "00"&x"0284E", "11"&x"FF756", "11"&x"FE261", "00"&x"02EB3", "11"&x"FE215", "11"&x"FF729", "00"&x"02989", "11"&x"FD3B6", "00"&x"00ECA", "00"&x"019C4", "11"&x"FD00F", 
                                "00"&x"02364", "00"&x"00310", "11"&x"FD85A", "00"&x"02FAF", "11"&x"FEAF0", "11"&x"FEAD8", "00"&x"03058", "11"&x"FD770", "00"&x"00329", "00"&x"024DF", "11"&x"FCD97", "00"&x"01B57", "00"&x"00FD6", "11"&x"FD024", "00"&x"02D4C", "11"&x"FF645", 
                                "11"&x"FDEC5", "00"&x"03458", "11"&x"FDE7E", "11"&x"FF61C", "00"&x"02E70", "11"&x"FCE86", "00"&x"01082", "00"&x"01CBD", "11"&x"FCA93", "00"&x"02768", "00"&x"00368", "11"&x"FD3EC", "00"&x"034F8", "11"&x"FE8A0", "11"&x"FE889", "00"&x"03593", 
                                "11"&x"FD315", "00"&x"0037F", "00"&x"028C4", "11"&x"FC84F", "00"&x"01E2F", "00"&x"01178", "11"&x"FCB3F", "00"&x"031E4", "11"&x"FF54B", "11"&x"FDB74", "00"&x"03987", "11"&x"FDB34", "11"&x"FF525", "00"&x"032EC", "11"&x"FC9C9", "00"&x"01213", 
                                "00"&x"01F72", "11"&x"FC595", "00"&x"02B0F", "00"&x"003B8", "11"&x"FCFE8", "00"&x"039C1", "11"&x"FE688", "11"&x"FE674", "00"&x"03A4A", "11"&x"FCF2A", "00"&x"003CD", "00"&x"02C44", "11"&x"FC393", "00"&x"020BA", "00"&x"012EE", "11"&x"FC6E0", 
                                "00"&x"035FD", "11"&x"FF46C", "11"&x"FD881", "00"&x"03E20", "11"&x"FD84A", "11"&x"FF44B", "00"&x"036E3", "11"&x"FC59B", "00"&x"01375", "00"&x"021D4", "11"&x"FC133", "00"&x"02E42", "00"&x"003FE", "11"&x"FCC66", "00"&x"03DEE", "11"&x"FE4B5", 
                                "11"&x"FE4A4", "00"&x"03E63", "11"&x"FCBC3", "00"&x"00410", "00"&x"02F4A", "11"&x"FBF7D", "00"&x"022EB", "00"&x"0142F", "11"&x"FC321", "00"&x"0397F", "11"&x"FF3AD", "11"&x"FD5FE", "00"&x"0420B", "11"&x"FD5CF", "11"&x"FF392", "00"&x"03A3E", 
                                "11"&x"FC213", "00"&x"0149F", "00"&x"023D4", "11"&x"FBD85", "00"&x"030F1", "00"&x"00439", "11"&x"FC979", "00"&x"04167", "11"&x"FE331", "11"&x"FE323", "00"&x"041C5", "11"&x"FC8F6", "00"&x"00447", "00"&x"031C4", "11"&x"FBC26", "00"&x"024B5", 
                                "00"&x"01534", "11"&x"FC016", "00"&x"03C56", "11"&x"FF313", "11"&x"FD3F7", "00"&x"04530", "11"&x"FD3D4", "11"&x"FF2FE", "00"&x"03CE9", "11"&x"FBF46", "00"&x"0158B", "00"&x"02569", "11"&x"FBAA1", "00"&x"0330A", "00"&x"00467", "11"&x"FC732", 
                                "00"&x"04419", "11"&x"FE206", "11"&x"FE1FC", "00"&x"0445D", "11"&x"FC6D3", "00"&x"00471", "00"&x"033A5", "11"&x"FB9A0", "00"&x"0260D", "00"&x"015F8", "11"&x"FBDD2", "00"&x"03E71", "11"&x"FF2A2", "11"&x"FD27B", "00"&x"0477C", "11"&x"FD262", 
                                "11"&x"FF293", "00"&x"03ED5", "11"&x"FBD44", "00"&x"01633", "00"&x"02687", "11"&x"FB898", "00"&x"03482", "00"&x"00486", "11"&x"FC59F", "00"&x"045F2", "11"&x"FE13A", "11"&x"FE134", "00"&x"0461B", "11"&x"FC565", "00"&x"0048D", "00"&x"034E0", 
                                "11"&x"FB7FC", "00"&x"026EB", "00"&x"01675", "11"&x"FBC61", "00"&x"03FC4", "11"&x"FF25B", "11"&x"FD190", "00"&x"048E2", "11"&x"FD184", "11"&x"FF254", "00"&x"03FF6", "11"&x"FBC1A", "00"&x"01693", "00"&x"02729", "11"&x"FB776", "00"&x"03550", 
                                "00"&x"00498", "11"&x"FC4CA", "00"&x"046E8", "11"&x"FE0D2", "11"&x"FE0CF", "00"&x"046F6", "11"&x"FC4B6", "00"&x"0049A", "00"&x"03570", "11"&x"FB742", "00"&x"0274A", "00"&x"016A9", "11"&x"FBBCE", "00"&x"04046", "11"&x"FF241", "11"&x"FD13D", 
                                "00"&x"0495B", "11"&x"FD13D", "11"&x"FF241", "00"&x"04046", "11"&x"FBBCE", "00"&x"016A9", "00"&x"0274A", "11"&x"FB742", "00"&x"03570", "00"&x"0049A", "11"&x"FC4B6", "00"&x"046F6", "11"&x"FE0CF", "11"&x"FE0D2", "00"&x"046E8", "11"&x"FC4CA", 
                                "00"&x"00498", "00"&x"03550", "11"&x"FB776", "00"&x"02729", "00"&x"01693", "11"&x"FBC1A", "00"&x"03FF6", "11"&x"FF254", "11"&x"FD184", "00"&x"048E2", "11"&x"FD190", "11"&x"FF25B", "00"&x"03FC4", "11"&x"FBC61", "00"&x"01675", "00"&x"026EB", 
                                "11"&x"FB7FC", "00"&x"034E0", "00"&x"0048D", "11"&x"FC565", "00"&x"0461B", "11"&x"FE134", "11"&x"FE13A", "00"&x"045F2", "11"&x"FC59F", "00"&x"00486", "00"&x"03482", "11"&x"FB898", "00"&x"02687", "00"&x"01633", "11"&x"FBD44", "00"&x"03ED5", 
                                "11"&x"FF293", "11"&x"FD262", "00"&x"0477C", "11"&x"FD27B", "11"&x"FF2A2", "00"&x"03E71", "11"&x"FBDD2", "00"&x"015F8", "00"&x"0260D", "11"&x"FB9A0", "00"&x"033A5", "00"&x"00471", "11"&x"FC6D3", "00"&x"0445D", "11"&x"FE1FC", "11"&x"FE206", 
                                "00"&x"04419", "11"&x"FC732", "00"&x"00467", "00"&x"0330A", "11"&x"FBAA1", "00"&x"02569", "00"&x"0158B", "11"&x"FBF46", "00"&x"03CE9", "11"&x"FF2FE", "11"&x"FD3D4", "00"&x"04530", "11"&x"FD3F7", "11"&x"FF313", "00"&x"03C56", "11"&x"FC016", 
                                "00"&x"01534", "00"&x"024B5", "11"&x"FBC26", "00"&x"031C4", "00"&x"00447", "11"&x"FC8F6", "00"&x"041C5", "11"&x"FE323", "11"&x"FE331", "00"&x"04167", "11"&x"FC979", "00"&x"00439", "00"&x"030F1", "11"&x"FBD85", "00"&x"023D4", "00"&x"0149F", 
                                "11"&x"FC213", "00"&x"03A3E", "11"&x"FF392", "11"&x"FD5CF", "00"&x"0420B", "11"&x"FD5FE", "11"&x"FF3AD", "00"&x"0397F", "11"&x"FC321", "00"&x"0142F", "00"&x"022EB", "11"&x"FBF7D", "00"&x"02F4A", "00"&x"00410", "11"&x"FCBC3", "00"&x"03E63", 
                                "11"&x"FE4A4", "11"&x"FE4B5", "00"&x"03DEE", "11"&x"FCC66", "00"&x"003FE", "00"&x"02E42", "11"&x"FC133", "00"&x"021D4", "00"&x"01375", "11"&x"FC59B", "00"&x"036E3", "11"&x"FF44B", "11"&x"FD84A", "00"&x"03E20", "11"&x"FD881", "11"&x"FF46C", 
                                "00"&x"035FD", "11"&x"FC6E0", "00"&x"012EE", "00"&x"020BA", "11"&x"FC393", "00"&x"02C44", "00"&x"003CD", "11"&x"FCF2A", "00"&x"03A4A", "11"&x"FE674", "11"&x"FE688", "00"&x"039C1", "11"&x"FCFE8", "00"&x"003B8", "00"&x"02B0F", "11"&x"FC595", 
                                "00"&x"01F72", "00"&x"01213", "11"&x"FC9C9", "00"&x"032EC", "11"&x"FF525", "11"&x"FDB34", "00"&x"03987", "11"&x"FDB74", "11"&x"FF54B", "00"&x"031E4", "11"&x"FCB3F", "00"&x"01178", "00"&x"01E2F", "11"&x"FC84F", "00"&x"028C4", "00"&x"0037F", 
                                "11"&x"FD315", "00"&x"03593", "11"&x"FE889", "11"&x"FE8A0", "00"&x"034F8", "11"&x"FD3EC", "00"&x"00368", "00"&x"02768", "11"&x"FCA93", "00"&x"01CBD", "00"&x"01082", "11"&x"FCE86", "00"&x"02E70", "11"&x"FF61C", "11"&x"FDE7E", "00"&x"03458", 
                                "11"&x"FDEC5", "11"&x"FF645", "00"&x"02D4C", "11"&x"FD024", "00"&x"00FD6", "00"&x"01B57", "11"&x"FCD97", "00"&x"024DF", "00"&x"00329", "11"&x"FD770", "00"&x"03058", "11"&x"FEAD8", "11"&x"FEAF0", "00"&x"02FAF", "11"&x"FD85A", "00"&x"00310", 
                                "00"&x"02364", "11"&x"FD00F", "00"&x"019C4", "00"&x"00ECA", "11"&x"FD3B6", "00"&x"02989", "11"&x"FF729", "11"&x"FE215", "00"&x"02EB3", "11"&x"FE261", "11"&x"FF756", "00"&x"0284E", "11"&x"FD573", "00"&x"00E11", "00"&x"01844", "11"&x"FD34D", 
                                "00"&x"020AB", "00"&x"002CC", "11"&x"FDC20", "00"&x"02AB7", "11"&x"FED53", "11"&x"FED6D", "00"&x"02A04", "11"&x"FDD19", "00"&x"002B1", "00"&x"01F18", "11"&x"FD5EA", "00"&x"01699", "00"&x"00CF5", "11"&x"FD93C", "00"&x"02451", "11"&x"FF847", 
                                "11"&x"FE5E4", "00"&x"028B6", "11"&x"FE634", "11"&x"FF876", "00"&x"02308", "11"&x"FDB0E", "00"&x"00C33", "00"&x"01506", "11"&x"FD950", "00"&x"01C3E", "00"&x"0026A", "11"&x"FE10D", "00"&x"024CF", "11"&x"FEFEC", "11"&x"FF007", "00"&x"02417", 
                                "11"&x"FE20E", "00"&x"0024E", "00"&x"01A9E", "11"&x"FDC05", "00"&x"0134C", "00"&x"00B0D", "11"&x"FDEFA", "00"&x"01EE7", "11"&x"FF970", "11"&x"FE9D6", "00"&x"02284", "11"&x"FEA28", "11"&x"FF9A0", "00"&x"01D96", "11"&x"FE0D6", "00"&x"00A47", 
                                "00"&x"011B0", "11"&x"FDF7F", "00"&x"017B2", "00"&x"00206", "11"&x"FE61A", "00"&x"01EC2", "11"&x"FF295", "11"&x"FF2B1", "00"&x"01E07", "11"&x"FE71F", "00"&x"001EA", "00"&x"0160C", "11"&x"FE23D", "00"&x"00FF0", "00"&x"0091D", "11"&x"FE4CF", 
                                "00"&x"01968", "11"&x"FFA9D", "11"&x"FEDD6", "00"&x"01C3D", "11"&x"FEE28", "11"&x"FFACD", "00"&x"01816", "11"&x"FE6AC", "00"&x"00856", "00"&x"00E53", "11"&x"FE5B8", "00"&x"01320", "00"&x"001A1", "11"&x"FEB2D", "00"&x"018AF", "11"&x"FF541", 
                                "11"&x"FF55C", "00"&x"017F6", "11"&x"FEC2F", "00"&x"00185", "00"&x"0117D", "11"&x"FE871", "00"&x"00C97", "00"&x"0072F", "11"&x"FEA9C", "00"&x"013F0", "11"&x"FFBC8", "11"&x"FF1CF", "00"&x"01603", "11"&x"FF21F", "11"&x"FFBF7", "00"&x"012A5", 
                                "11"&x"FEC71", "00"&x"0066C", "00"&x"00B01", "11"&x"FEBDC", "00"&x"00E9E", "00"&x"0013E", "11"&x"FF02B", "00"&x"012B7", "11"&x"FF7E0", "11"&x"FF7FA", "00"&x"01203", "11"&x"FF126", "00"&x"00123", "00"&x"00D07", "11"&x"FEE80", "00"&x"00952", 
                                "00"&x"0054D", "11"&x"FF045", "00"&x"00E9D", "11"&x"FFCEB", "11"&x"FF5AB", "00"&x"00FF7", "11"&x"FF5F9", "11"&x"FFD18", "00"&x"00D5E", "11"&x"FF208", "00"&x"00491", "00"&x"007CC", "11"&x"FF1CA", "00"&x"00A44", "00"&x"000DE", "11"&x"FF4FA", 
                                "00"&x"00CF8", "11"&x"FFA65", "11"&x"FFA7E", "00"&x"00C4D", "11"&x"FF5E9", "00"&x"000C4", "00"&x"008C2", "11"&x"FF44E", "00"&x"00631", "00"&x"00380", "11"&x"FF5AB", "00"&x"00989", "11"&x"FFE00", "11"&x"FF959", "00"&x"00A36", "11"&x"FF9A1", 
                                "11"&x"FFE2B", "00"&x"0085D", "11"&x"FF754", "00"&x"002D0", "00"&x"004C3", "11"&x"FF766", "00"&x"00629", "00"&x"00084", "11"&x"FF983", "00"&x"0078E", "11"&x"FFCC5", "11"&x"FFCDC", "00"&x"006EF", "11"&x"FFA61", "00"&x"0006C", "00"&x"004C1", 
                                "11"&x"FF9BC", "00"&x"00345", "00"&x"001D2", "11"&x"FFAB6", "00"&x"004CC", "11"&x"FFF03", "11"&x"FFCC5", "00"&x"004DB", "11"&x"FFD08", "11"&x"FFF2A", "00"&x"003B9", "11"&x"FFC3C", "00"&x"00130", "00"&x"001F3", "11"&x"FFC95", "00"&x"0025D", 
                                "00"&x"00031", "11"&x"FFDB1", "00"&x"00292", "11"&x"FFEF3", "11"&x"FFF09", "00"&x"00201", "11"&x"FFE7A", "00"&x"0001B", "00"&x"00117", "11"&x"FFEB4", "00"&x"00099", "00"&x"00049", "11"&x"FFF4F", "00"&x"0007C", "11"&x"FFFEE", "11"&x"FFFE1", 
                                "11"&x"FFFFF", "00"&x"0001D", "00"&x"00011", "11"&x"FFF85", "00"&x"000AC", "11"&x"FFFB8", "11"&x"FFF6B", "00"&x"00140", "11"&x"FFEF3", "11"&x"FFFE6", "00"&x"00172", "11"&x"FFE19", "00"&x"000E8", "00"&x"000FB", "11"&x"FFD9A", "00"&x"00223", 
                                "11"&x"FFFD2", "11"&x"FFDD3", "00"&x"0031F", "11"&x"FFE39", "11"&x"FFEEC", "00"&x"00363", "11"&x"FFCAA", "00"&x"000BE", "00"&x"002A1", "11"&x"FFBB6", "00"&x"002D5", "00"&x"000DC", "11"&x"FFBD4", "00"&x"00492", "11"&x"FFE6E", "11"&x"FFD33", 
                                "00"&x"00555", "11"&x"FFBF8", "11"&x"FFFA4", "00"&x"004B7", "11"&x"FFA36", "00"&x"0029B", "00"&x"002AB", "11"&x"FF9C9", "00"&x"0054E", "11"&x"FFF94", "11"&x"FFB02", "00"&x"006EE", "11"&x"FFC2E", "11"&x"FFDC1", "00"&x"006E1", "11"&x"FF964", 
                                "00"&x"00170", "00"&x"004FA", "11"&x"FF80E", "00"&x"00525", "00"&x"00189", "11"&x"FF8B1", "00"&x"007DF", "11"&x"FFD58", "11"&x"FFB53", "00"&x"008C6", "11"&x"FF975", "11"&x"FFF6D", "00"&x"00775", "11"&x"FF6F4", "00"&x"00407", "00"&x"00414", 
                                "11"&x"FF69B", "00"&x"007F0", "11"&x"FFF60", "11"&x"FF8AD", "00"&x"00A14", "11"&x"FFA7E", "11"&x"FFCCA", "00"&x"009C1", "11"&x"FF6B5", "00"&x"00201", "00"&x"006E5", "11"&x"FF513", "00"&x"00707", "00"&x"00216", "11"&x"FF627", "00"&x"00A8A", 
                                "11"&x"FFC77", "11"&x"FF9D1", "00"&x"00B8B", "11"&x"FF772", "11"&x"FFF41", "00"&x"009A5", "11"&x"FF45C", "00"&x"00527", "00"&x"00531", "11"&x"FF418", "00"&x"00A03", "11"&x"FFF37", "11"&x"FF6D9", "00"&x"00C8A", "11"&x"FF92E", "11"&x"FFC0A", 
                                "00"&x"00BFC", "11"&x"FF4A1", "00"&x"00272", "00"&x"0085E", "11"&x"FF2CA", "00"&x"00877", "00"&x"00280", "11"&x"FF439", "00"&x"00C8F", "11"&x"FFBCD", "11"&x"FF8AF", "00"&x"00D9D", "11"&x"FF5F2", "11"&x"FFF21", "00"&x"00B44", "11"&x"FF272"
    );

    -- 24 bit accumulator
    signal accumulator : sfixed(0 downto -23) := (others => '0');
    -- 12 bit because max sum is 1286.28
    --signal accumulator : signed(23 downto 0) := (others => '0');
    signal sfixed_data_in : sfixed(0 downto 0) := (others => '0');

    signal tap_counter : unsigned(11 downto 0) := (others => '0');
    

begin

    FIR_PROC : process(clk)

        variable v_prev_ready : std_logic := '0';
        variable v_next_valid : std_logic := '0';
        variable v_index : integer range 0 to FIR_LENGTH * 2 - 1 := 0;
        variable v_coeff : sfixed(0 downto -21);
        variable v_delay_line : sfixed(0 downto 0);
        variable v_mult_result : sfixed(0 downto -21);

    begin
        
        if rising_edge(clk) then

            -- Default values
            v_prev_ready := '0';
            v_next_valid := '0';

            if rst_n = '0' then

                state <= IDLE;
                
            else
                
                case state is

                    -------------------------------
                    when IDLE =>
                        -------------------------------
                        v_prev_ready := '1';

                        if prev_valid = '1' then
                            state <= SHIFT_DATA_IN;
                        end if;

                    -------------------------------
                    when SHIFT_DATA_IN =>
                        -------------------------------
                        delay_line <= data_in & delay_line(delay_line'low to delay_line'high - 1);

                        -- Get accumulator ready
                        accumulator <=  (others => '0');
                        state <= CALCULATE;


                    -------------------------------
                    when CALCULATE =>
                        -------------------------------

                        v_index := to_integer(tap_counter);

                        v_coeff := coeff(v_index);
                        v_delay_line := to_sfixed(delay_line(v_index)(0 downto 0), v_delay_line);

                        v_mult_result := resize(v_coeff * v_delay_line , v_mult_result); -- * to_sfixed(-1, v_delay_line)

                        accumulator <= resize(accumulator + v_mult_result, accumulator);--fixed_saturate, fixed_round);

                        if (tap_counter < FIR_LENGTH - 1) then
                            tap_counter <= tap_counter + 1;
                        else
                            tap_counter <= (others => '0');
                            state <= HOLD_DATA_OUT;
                        end if;

                    -------------------------------
                    when HOLD_DATA_OUT =>
                        -------------------------------
                        v_next_valid := '1';

                        data_out <= accumulator;
                        
                        if next_ready = '1' then
                            state <= IDLE;
                        end if;

                end case;

            end if;

            prev_ready <= v_prev_ready;
            next_valid <= v_next_valid;

        end if;
        
    end process;

end architecture;